package tb_decryptor_pkg;
    import uvm_pkg::*;
`include "uvm_macros.svh"
`include "tb_ip_item.svh"
`include "tb_op_item.svh"
`include "tb_cfg_item.svh"
`include "tb_var_len_item.svh"
`include "tb_var_init_item.svh"

`include "def_sequence.svh"
`include "tb_mem_test_seq.svh"
`include "tb_rand_seq.svh"

`include "tb_driver_uvm.svh"
`include "tb_monitor_uvm.svh"
`include "tb_scoreboard_uvm.svh"
`include "coverage.svh"

`include "tb_env_uvm.svh"

`include "tb_base_test.svh"
`include "tb_smoketest.svh"
`include "tb_mem_test.svh"
`include "tb_rand_test.svh"
`include "tb_var_len_test.svh"
`include "tb_var_init_test.svh"
`include "tb_parallel_test.svh"
endpackage